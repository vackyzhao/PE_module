module fpga_top (
    input clk,
    input rst_n,
    input i_cam
);
    
endmodule