module PingPongBuffer();

endmodule 