//Copyright (C)2014-2022 Gowin Semiconductor Corporation.
//All rights reserved.
//File Title: IP file
//GOWIN Version: V1.9.8.07 Education
//Part Number: GW2A-LV18PG256C8/I7
//Device: GW2A-18C
//Created Time: Thu Aug 18 22:10:45 2022

module cmos_pll (clkout, clkin);

output clkout;
input clkin;

assign clkout=clkin;

endmodule //cmos_pll
